module uart(
  
)
endmodule